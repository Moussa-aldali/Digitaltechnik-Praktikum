library ieee;
use ieee.std_logic_1164.all;

entity zeiger is
  port(
     x: in std_logic_vector (4 downto 0);
     segments: out std_logic_vector (6 downto 0));
 end zeiger;
 
architecture arch of zeiger is
begin
 with x select ---------------------------0--------------------------------- 
  segments <= "0000001" when "00000",
              ---------------------------1---------------------------------- 
              "1001111" when "00001",
              ---------------------------2---------------------------------- 
              "0010010" when "00010",
              ---------------------------3---------------------------------- 
              "0000110" when "00011",
              ---------------------------4---------------------------------- 
              "1001100" when "00100",
              ---------------------------5---------------------------------- 
              "0100100" when "00101",
              ---------------------------6---------------------------------- 
              "0100000" when "00110",
              ---------------------------7---------------------------------- 
              "0001101" when "00111",
              ---------------------------8---------------------------------- 
              "0000000" when "01000",
              ---------------------------9---------------------------------- 
              "0000100" when "01001",
              ---------------------------10---------------------------------- P
              "0011000" when "01010",
              ---------------------------11---------------------------------- N
              "0001001" when "01011",
              ---------------------------12---------------------------------- C
              "0110001" when "01100",
              ---------------------------13----------------------------------  D
              "1000010" when "01101",
              ---------------------------14----------------------------------  E
              "0110000" when "01110",
              ---------------------------15---------------------------------- R
              "1111010" when "01111",
              ---------------------------16---------------------------------- L
              "1110001" when "10000",
              ---------------------------17----------------------------------  BLANKEN
              "0110110" when "10001",
              ---------------------------18---------------------------------- 
              "1111111" when others;
            
end arch;

